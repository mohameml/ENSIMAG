library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity FD8CE is
    port (
        Q   : out unsigned(7 downto 0) := (others => '0');
        C   : in STD_LOGIC;
        CE  : in STD_LOGIC;
        CLR : in STD_LOGIC;
        D   : in unsigned(7 downto 0)
    );
end FD8CE;

architecture Behavioral of FD8CE is
begin
    process(C, CLR)
    begin
        if (CLR='1') then
            Q <= (others => '0');
        elsif (C'event and C = '1') then
            if (CE='1') then
                Q <= D;
            end if;
        end if;
    end process;
end Behavioral;
